C:\TRANSFER\tmp4\IBIST1.cir Setup1
*#save V(400) @V4[i] @V4[p] V(100) @V1[i] @V1[p] V(500) @V2[i]
*#save @V2[p] V(7) @C1[i] @C1[p] V(300) @V3[i] @V3[p]
*#alias vpcebb  v(7)
*#VIEW  TRAN vpcebb
*#alias V_100  v(100)
*#VIEW  TRAN V_100
*#alias V_500  v(500)
*#VIEW  TRAN V_500
.TRAN .1n 120n 0 1n UIC
.OPTIONS itl1=300
.PRINT  TRAN vpcebb
.PRINT  TRAN V_100
.PRINT  TRAN V_500
V4 400 0 DC=0
V1 100 0 PULSE 0 5 0 2.5N 2.5N 27.44N 59.88N 
V2 500 0 DC=5
C1 7 0 50PF
V3 300 0 DC=5
X4 100 7 300 400 500 PCEBB12211_W {  }
.SUBCKT PCEBB12211_W 100 4 300 400 500
*Connections    Input Output VCC VEE Enable
;
; E:\SPICE4\CIRCUITS\APPS\IBIS\82375sb.ibs
; Tuesday, September 08, 1998 15:33:41
;
; Referenced by:
; LA31, LA30, LA29, LA28, LA27
; LA26, LA25, LA24, LA16, LA15
; LA14, LA13, LA12, LA11, LA10
; LA9, LA8, LA7, LA6, LA5
; LA4, LA23, LA3, LA22, LA2
; LA21, LA20, LA19, LA18, LA17
; AD31, AD30, AD29, AD28, AD27
; AD26, AD25, AD24, C/BE3#, AD23
; AD22, AD21, AD20, AD19, AD18
; AD17, AD16, C/BE2#, FRAME#, IRDY#
; TRDY#, DEVSEL#, STOP#, PCILOCK#, PERR#
; PAR, C/BE1#, AD15, AD14, AD13
; AD12, AD11, AD10, AD9, C/BE0#
; AD8, AD7, AD6, AD5, AD4
; AD3, AD2, AD1, AD0, LOCK#
; START#, EXRDY, SLBURST#, MSBURST#, M/IO#
; W/R#, BE3#, BE2#, BE1#, BE0#
*Passed Parameters; worst
*DEFINE {RTF}=  30.079k  ;2.84V/854.23ps
*DEFINE {RTR}=  23.849k  ;2.27V/541.37ps
* Input Control
B1 820 0 V=V(100) & V(500)
B2 830 0 V= V(500) & ~V(100)
* Up and Down Ramps
B3 300 850 I= V(830) > 1.2   ? 0 : V(300,850) / {RTR}
B4 840 400 I= V(820) > 1.2 ? 0 : V(840,400) / {RTF}
C1 300 850 .01P
C2 840 400 .01P
S1 220 850 0 820 SMOD
S2 840 220 0 830 SMOD
.MODEL SMOD SW RON=.1M ROFF=1E15 VT=-1.2 VH=.1
G1 8 400 2 8 1
R1 6 400 1
G2 300 8 8 3 1
R2 300 6 1
* Pull-up/Pull-down structures; worst

XEPL_DN 2 400 8 840 PULL_DOWN


XEPL_UP 3 300 850 8 PULL_UP

* Diode Clamps

XPWR_CLAMP 6 300 300 6 PWR_CLAMP


XGND_OUT 6 400 6 400 GND_CLAMP

* Package Parasitics; worst
ROSNB 5 1 100
ROPKG 1 4 277.0m
COPKG 4 400 2.11pF
CCOMP 5 400 4.28pF
LOPKG 5 1 14.76nH
* Voltage Sources for measuring currents
V5 6 5 
V6 8 6 
V7 220 8 
.ENDS


.SUBCKT	GND_CLAMP	3    4   1   2
; connections:      Out+ Out In+ In
B1	3 4	I=
+ (V(1,2) <   -5.000 ) ?    1.000n * V(1,2) +  -84.800  : 
+ (V(1,2) <   -4.800 ) ?   20.900  * V(1,2) +   19.700  : 
+ (V(1,2) <   -4.600 ) ?   20.850  * V(1,2) +   19.460  : 
+ (V(1,2) <   -4.400 ) ?   20.900  * V(1,2) +   19.690  : 
+ (V(1,2) <   -4.200 ) ?   20.850  * V(1,2) +   19.470  : 
+ (V(1,2) <   -4.000 ) ?   20.850  * V(1,2) +   19.470  : 
+ (V(1,2) <   -3.800 ) ?   20.800  * V(1,2) +   19.270  : 
+ (V(1,2) <   -3.600 ) ?   20.850  * V(1,2) +   19.460  : 
+ (V(1,2) <   -3.400 ) ?   20.800  * V(1,2) +   19.280  : 
+ (V(1,2) <   -3.200 ) ?   20.800  * V(1,2) +   19.280  : 
+ (V(1,2) <   -3.000 ) ?   20.750  * V(1,2) +   19.120  : 
+ (V(1,2) <   -2.800 ) ?   20.750  * V(1,2) +   19.120  : 
+ (V(1,2) <   -2.600 ) ?   20.700  * V(1,2) +   18.980  : 
+ (V(1,2) <   -2.400 ) ?   20.700  * V(1,2) +   18.980  : 
+ (V(1,2) <   -2.200 ) ?   20.650  * V(1,2) +   18.860  : 
+ (V(1,2) <   -2.000 ) ?   20.600  * V(1,2) +   18.750  : 
+ (V(1,2) <   -1.950 ) ?   20.400  * V(1,2) +   18.350  : 
+ (V(1,2) <   -1.900 ) ?   20.600  * V(1,2) +   18.740  : 
+ (V(1,2) <   -1.850 ) ?   20.400  * V(1,2) +   18.360  : 
+ (V(1,2) <   -1.800 ) ?   20.600  * V(1,2) +   18.730  : 
+ (V(1,2) <   -1.750 ) ?   20.400  * V(1,2) +   18.370  : 
+ (V(1,2) <   -1.700 ) ?   20.400  * V(1,2) +   18.370  : 
+ (V(1,2) <   -1.650 ) ?   20.400  * V(1,2) +   18.370  : 
+ (V(1,2) <   -1.600 ) ?   20.200  * V(1,2) +   18.040  : 
+ (V(1,2) <   -1.550 ) ?   20.400  * V(1,2) +   18.360  : 
+ (V(1,2) <   -1.500 ) ?   20.200  * V(1,2) +   18.050  : 
+ (V(1,2) <   -1.450 ) ?   20.000  * V(1,2) +   17.750  : 
+ (V(1,2) <   -1.400 ) ?   20.200  * V(1,2) +   18.040  : 
+ (V(1,2) <   -1.350 ) ?   20.000  * V(1,2) +   17.760  : 
+ (V(1,2) <   -1.300 ) ?   19.800  * V(1,2) +   17.490  : 
+ (V(1,2) <   -1.250 ) ?   19.800  * V(1,2) +   17.490  : 
+ (V(1,2) <   -1.200 ) ?   19.600  * V(1,2) +   17.240  : 
+ (V(1,2) <   -1.150 ) ?   19.200  * V(1,2) +   16.760  : 
+ (V(1,2) <   -1.100 ) ?   19.200  * V(1,2) +   16.760  : 
+ (V(1,2) <   -1.050 ) ?   18.200  * V(1,2) +   15.660  : 
+ (V(1,2) <   -1.000 ) ?   18.400  * V(1,2) +   15.870  : 
+ (V(1,2) < -950.000m) ?   16.000  * V(1,2) +   13.470  : 
+ (V(1,2) < -900.000m) ?   16.050  * V(1,2) +   13.518  : 
+ (V(1,2) < -850.000m) ?    8.530  * V(1,2) +    6.750  : 
+ (V(1,2) < -800.000m) ?    8.530  * V(1,2) +    6.750  : 
+ (V(1,2) < -750.000m) ?  732.400m * V(1,2) +  511.450m : 
+ (V(1,2) < -700.000m) ?  732.200m * V(1,2) +  511.300m : 
+ (V(1,2) < -650.000m) ?   12.207m * V(1,2) +    7.305m : 
+ (V(1,2) < -600.000m) ?   12.225m * V(1,2) +    7.316m : 
+ (V(1,2) < -550.000m) ?  181.200u * V(1,2) +   90.290u : 
+ (V(1,2) < -500.000m) ?  181.122u * V(1,2) +   90.247u : 
+ (V(1,2) < -450.000m) ?    3.061u * V(1,2) +    1.217u : 
+ (V(1,2) < -400.000m) ?    3.061u * V(1,2) +    1.217u : 
+ (V(1,2) < -350.000m) ?   76.000n * V(1,2) +   22.600n : 
+ (V(1,2) < -300.000m) ?   75.940n * V(1,2) +   22.579n : 
+ (V(1,2) < -250.000m) ?    2.725n * V(1,2) +  614.380p : 
+ (V(1,2) < -200.000m) ?    2.725n * V(1,2) +  614.430p : 
+ (V(1,2) < -150.000m) ?  260.400p * V(1,2) +  121.550p : 
+ (V(1,2) < -100.000m) ?  260.600p * V(1,2) +  121.580p : 
+ (V(1,2) <  -50.000m) ? -197.600p * V(1,2) +   75.760p : 
+ (V(1,2) <    0.000 ) ? -197.600p * V(1,2) +   75.760p : 
+ (V(1,2) <    5.000 ) ?    5.060p * V(1,2) +   75.760p : 
+    1.000n * V(1,2) +  101.060p
.ENDS


.SUBCKT	PULL_UP	3    4   1   2
; connections:  Out+ Out In+ In
B1	3 4	V=
+ (V(1,2) <   -5.000 ) ?    1.000n * V(1,2) +  363.790u : 
+ (V(1,2) <   -4.500 ) ?   98.320u * V(1,2) +  855.390u : 
+ (V(1,2) <   -4.000 ) ?  129.360u * V(1,2) +  995.070u : 
+ (V(1,2) <   -3.500 ) ?  177.900u * V(1,2) +    1.189m : 
+ (V(1,2) <   -3.000 ) ?  260.100u * V(1,2) +    1.477m : 
+ (V(1,2) <   -2.500 ) ?  416.400u * V(1,2) +    1.946m : 
+ (V(1,2) <   -2.000 ) ?  770.340u * V(1,2) +    2.831m : 
+ (V(1,2) <   -1.500 ) ?    1.940m * V(1,2) +    5.170m : 
+ (V(1,2) <   -1.400 ) ?    3.900m * V(1,2) +    8.110m : 
+ (V(1,2) <   -1.300 ) ?    5.500m * V(1,2) +   10.350m : 
+ (V(1,2) <   -1.200 ) ?    8.600m * V(1,2) +   14.380m : 
+ (V(1,2) <   -1.100 ) ?   14.200m * V(1,2) +   21.100m : 
+ (V(1,2) <   -1.000 ) ?   28.500m * V(1,2) +   36.830m : 
+ (V(1,2) < -900.000m) ?   75.500m * V(1,2) +   83.830m : 
+ (V(1,2) < -800.000m) ?  238.700m * V(1,2) +  230.710m : 
+ (V(1,2) < -700.000m) ?   73.600m * V(1,2) +   98.630m : 
+ (V(1,2) < -600.000m) ?  -63.600m * V(1,2) +    2.590m : 
+ (V(1,2) < -500.000m) ?  -67.400m * V(1,2) +  310.000u : 
+ (V(1,2) < -400.000m) ?  -67.700m * V(1,2) +  160.000u : 
+ (V(1,2) < -300.000m) ?  -68.000m * V(1,2) +   40.000u : 
+ (V(1,2) < -200.000m) ?  -68.100m * V(1,2) +   10.000u : 
+ (V(1,2) < -100.000m) ?  -68.200m * V(1,2) +  -10.000u : 
+ (V(1,2) <    0.000 ) ?  -68.100m * V(1,2) +   -9.810p : 
+ (V(1,2) <  100.000m) ?  -67.100m * V(1,2) +   -9.810p : 
+ (V(1,2) <  200.000m) ?  -65.300m * V(1,2) + -180.000u : 
+ (V(1,2) <  300.000m) ?  -63.400m * V(1,2) + -560.000u : 
+ (V(1,2) <  400.000m) ?  -61.500m * V(1,2) +   -1.130m : 
+ (V(1,2) <  500.000m) ?  -59.700m * V(1,2) +   -1.850m : 
+ (V(1,2) <  600.000m) ?  -57.800m * V(1,2) +   -2.800m : 
+ (V(1,2) <  700.000m) ?  -56.000m * V(1,2) +   -3.880m : 
+ (V(1,2) <  800.000m) ?  -54.100m * V(1,2) +   -5.210m : 
+ (V(1,2) <  900.000m) ?  -52.200m * V(1,2) +   -6.730m : 
+ (V(1,2) <    1.000 ) ?  -50.400m * V(1,2) +   -8.350m : 
+ (V(1,2) <    1.100 ) ?  -48.500m * V(1,2) +  -10.250m : 
+ (V(1,2) <    1.200 ) ?  -46.600m * V(1,2) +  -12.340m : 
+ (V(1,2) <    1.300 ) ?  -44.800m * V(1,2) +  -14.500m : 
+ (V(1,2) <    1.400 ) ?  -42.900m * V(1,2) +  -16.970m : 
+ (V(1,2) <    1.500 ) ?  -41.000m * V(1,2) +  -19.630m : 
+ (V(1,2) <    1.600 ) ?  -39.200m * V(1,2) +  -22.330m : 
+ (V(1,2) <    1.700 ) ?  -37.300m * V(1,2) +  -25.370m : 
+ (V(1,2) <    1.800 ) ?  -35.300m * V(1,2) +  -28.770m : 
+ (V(1,2) <    1.900 ) ?  -33.600m * V(1,2) +  -31.830m : 
+ (V(1,2) <    2.000 ) ?  -31.700m * V(1,2) +  -35.440m : 
+ (V(1,2) <    2.100 ) ?  -29.800m * V(1,2) +  -39.240m : 
+ (V(1,2) <    2.200 ) ?  -28.000m * V(1,2) +  -43.020m : 
+ (V(1,2) <    2.300 ) ?  -26.100m * V(1,2) +  -47.200m : 
+ (V(1,2) <    2.400 ) ?  -24.300m * V(1,2) +  -51.340m : 
+ (V(1,2) <    2.500 ) ?  -22.400m * V(1,2) +  -55.900m : 
+ (V(1,2) <    2.600 ) ?  -20.500m * V(1,2) +  -60.650m : 
+ (V(1,2) <    2.700 ) ?  -18.600m * V(1,2) +  -65.590m : 
+ (V(1,2) <    2.800 ) ?  -16.800m * V(1,2) +  -70.450m : 
+ (V(1,2) <    2.900 ) ?  -15.000m * V(1,2) +  -75.490m : 
+ (V(1,2) <    3.000 ) ?  -13.000m * V(1,2) +  -81.290m : 
+ (V(1,2) <    3.100 ) ?  -11.200m * V(1,2) +  -86.690m : 
+ (V(1,2) <    3.200 ) ?   -9.300m * V(1,2) +  -92.580m : 
+ (V(1,2) <    3.300 ) ?   -7.500m * V(1,2) +  -98.340m : 
+ (V(1,2) <    3.400 ) ?   -5.600m * V(1,2) + -104.610m : 
+ (V(1,2) <    3.500 ) ?   -3.700m * V(1,2) + -111.070m : 
+ (V(1,2) <    3.600 ) ?  -11.400m * V(1,2) +  -84.120m : 
+ (V(1,2) <    3.700 ) ?  -14.500m * V(1,2) +  -72.960m : 
+ (V(1,2) <    3.800 ) ?   -9.400m * V(1,2) +  -91.830m : 
+ (V(1,2) <    3.900 ) ?   -7.900m * V(1,2) +  -97.530m : 
+ (V(1,2) <    4.000 ) ?   -7.000m * V(1,2) + -101.040m : 
+ (V(1,2) <    4.100 ) ?   -6.400m * V(1,2) + -103.440m : 
+ (V(1,2) <    4.200 ) ?   -5.900m * V(1,2) + -105.490m : 
+ (V(1,2) <    4.300 ) ?   -5.700m * V(1,2) + -106.330m : 
+ (V(1,2) <    4.400 ) ?   -5.400m * V(1,2) + -107.620m : 
+ (V(1,2) <    4.500 ) ?   -5.200m * V(1,2) + -108.500m : 
+ (V(1,2) <    4.600 ) ?   -5.000m * V(1,2) + -109.400m : 
+ (V(1,2) <    4.700 ) ?   -4.800m * V(1,2) + -110.320m : 
+ (V(1,2) <    4.800 ) ?   -4.800m * V(1,2) + -110.320m : 
+ (V(1,2) <    4.900 ) ?   -4.600m * V(1,2) + -111.280m : 
+ (V(1,2) <    5.000 ) ?   -4.600m * V(1,2) + -111.280m : 
+ (V(1,2) <    5.100 ) ?   -4.400m * V(1,2) + -112.280m : 
+ (V(1,2) <    5.200 ) ?   -4.400m * V(1,2) + -112.280m : 
+ (V(1,2) <    5.300 ) ?   -4.300m * V(1,2) + -112.800m : 
+ (V(1,2) <    5.400 ) ?   -4.200m * V(1,2) + -113.330m : 
+ (V(1,2) <    5.500 ) ?   -4.200m * V(1,2) + -113.330m : 
+ (V(1,2) <    5.600 ) ?   -4.100m * V(1,2) + -113.880m : 
+ (V(1,2) <    5.700 ) ?   -4.000m * V(1,2) + -114.440m : 
+ (V(1,2) <    5.800 ) ?   -4.100m * V(1,2) + -113.870m : 
+ (V(1,2) <    5.900 ) ?   -6.400m * V(1,2) + -100.530m : 
+ (V(1,2) <    6.000 ) ?  -89.500m * V(1,2) +  389.760m : 
+ (V(1,2) <    6.100 ) ?  355.800m * V(1,2) +   -2.282  : 
+ (V(1,2) <    6.200 ) ? -157.100m * V(1,2) +  846.650m : 
+ (V(1,2) <    6.300 ) ?  -87.900m * V(1,2) +  417.610m : 
+ (V(1,2) <    6.400 ) ?  -23.500m * V(1,2) +   11.890m : 
+ (V(1,2) <    6.500 ) ?  -12.100m * V(1,2) +  -61.070m : 
+ (V(1,2) <    7.000 ) ?   -4.620m * V(1,2) + -109.690m : 
+ (V(1,2) <    7.500 ) ?   -3.840m * V(1,2) + -115.150m : 
+ (V(1,2) <    8.000 ) ?   -3.580m * V(1,2) + -117.100m : 
+ (V(1,2) <    8.500 ) ?   -3.480m * V(1,2) + -117.900m : 
+ (V(1,2) <    9.000 ) ?   -3.420m * V(1,2) + -118.410m : 
+ (V(1,2) <    9.500 ) ?   -3.360m * V(1,2) + -118.950m : 
+ (V(1,2) <   10.000 ) ?   -3.260m * V(1,2) + -119.900m : 
+    1.000n * V(1,2) + -152.500m
.ENDS


.SUBCKT	PULL_DOWN	3    4   1   2
; connections:      Out+ Out In+ In
B1	3 4	V=
+ (V(1,2) <   -5.000 ) ?    1.000n * V(1,2) +   -1.060m : 
+ (V(1,2) <   -4.500 ) ? -300.000u * V(1,2) +   -2.560m : 
+ (V(1,2) <   -4.000 ) ? -380.000u * V(1,2) +   -2.920m : 
+ (V(1,2) <   -3.500 ) ? -520.000u * V(1,2) +   -3.480m : 
+ (V(1,2) <   -3.000 ) ? -780.000u * V(1,2) +   -4.390m : 
+ (V(1,2) <   -2.500 ) ?   -1.260m * V(1,2) +   -5.830m : 
+ (V(1,2) <   -2.000 ) ?   -2.360m * V(1,2) +   -8.580m : 
+ (V(1,2) <   -1.500 ) ?   -6.080m * V(1,2) +  -16.020m : 
+ (V(1,2) <   -1.400 ) ?  -12.700m * V(1,2) +  -25.950m : 
+ (V(1,2) <   -1.300 ) ?  -18.200m * V(1,2) +  -33.650m : 
+ (V(1,2) <   -1.200 ) ?  -28.900m * V(1,2) +  -47.560m : 
+ (V(1,2) <   -1.100 ) ?  -50.400m * V(1,2) +  -73.360m : 
+ (V(1,2) <   -1.000 ) ? -107.400m * V(1,2) + -136.060m : 
+ (V(1,2) < -900.000m) ? -319.000m * V(1,2) + -347.660m : 
+ (V(1,2) < -800.000m) ? -784.900m * V(1,2) + -766.970m : 
+ (V(1,2) < -700.000m) ?  -14.300m * V(1,2) + -150.490m : 
+ (V(1,2) < -600.000m) ?  173.900m * V(1,2) +  -18.750m : 
+ (V(1,2) < -500.000m) ?  184.400m * V(1,2) +  -12.450m : 
+ (V(1,2) < -400.000m) ?  192.200m * V(1,2) +   -8.550m : 
+ (V(1,2) < -300.000m) ?  200.300m * V(1,2) +   -5.310m : 
+ (V(1,2) < -200.000m) ?  208.700m * V(1,2) +   -2.790m : 
+ (V(1,2) < -100.000m) ?  217.900m * V(1,2) + -950.000u : 
+ (V(1,2) <    0.000 ) ?  227.400m * V(1,2) +    7.100n : 
+ (V(1,2) <  100.000m) ?  224.900m * V(1,2) +    7.100n : 
+ (V(1,2) <  200.000m) ?  210.300m * V(1,2) +    1.460m : 
+ (V(1,2) <  300.000m) ?  196.300m * V(1,2) +    4.260m : 
+ (V(1,2) <  400.000m) ?  183.100m * V(1,2) +    8.220m : 
+ (V(1,2) <  500.000m) ?  170.500m * V(1,2) +   13.260m : 
+ (V(1,2) <  600.000m) ?  158.600m * V(1,2) +   19.210m : 
+ (V(1,2) <  700.000m) ?  147.000m * V(1,2) +   26.170m : 
+ (V(1,2) <  800.000m) ?  136.200m * V(1,2) +   33.730m : 
+ (V(1,2) <  900.000m) ?  125.800m * V(1,2) +   42.050m : 
+ (V(1,2) <    1.000 ) ?  115.800m * V(1,2) +   51.050m : 
+ (V(1,2) <    1.100 ) ?  106.300m * V(1,2) +   60.550m : 
+ (V(1,2) <    1.200 ) ?   97.300m * V(1,2) +   70.450m : 
+ (V(1,2) <    1.300 ) ?   88.600m * V(1,2) +   80.890m : 
+ (V(1,2) <    1.400 ) ?   80.300m * V(1,2) +   91.680m : 
+ (V(1,2) <    1.500 ) ?   72.300m * V(1,2) +  102.880m : 
+ (V(1,2) <    1.600 ) ?   64.700m * V(1,2) +  114.280m : 
+ (V(1,2) <    1.700 ) ?   57.300m * V(1,2) +  126.120m : 
+ (V(1,2) <    1.800 ) ?   49.900m * V(1,2) +  138.700m : 
+ (V(1,2) <    1.900 ) ?   43.700m * V(1,2) +  149.860m : 
+ (V(1,2) <    2.000 ) ?   37.200m * V(1,2) +  162.210m : 
+ (V(1,2) <    2.100 ) ?   31.100m * V(1,2) +  174.410m : 
+ (V(1,2) <    2.200 ) ?   25.100m * V(1,2) +  187.010m : 
+ (V(1,2) <    2.300 ) ?   19.400m * V(1,2) +  199.550m : 
+ (V(1,2) <    2.400 ) ?    7.000m * V(1,2) +  228.070m : 
+ (V(1,2) <    2.500 ) ?    2.100m * V(1,2) +  239.830m : 
+ (V(1,2) <    2.600 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    2.700 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    2.800 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    2.900 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.000 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.100 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.200 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.300 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.400 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.500 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.600 ) ?    1.800m * V(1,2) +  240.580m : 
+ (V(1,2) <    3.700 ) ?    1.700m * V(1,2) +  240.940m : 
+ (V(1,2) <    3.800 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    3.900 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.000 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.100 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.200 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.300 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.400 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.500 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.600 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.700 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.800 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    4.900 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    5.000 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    5.100 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    5.200 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    5.300 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    5.400 ) ?    1.800m * V(1,2) +  240.570m : 
+ (V(1,2) <    5.500 ) ?    1.700m * V(1,2) +  241.110m : 
+ (V(1,2) <    5.600 ) ?    1.800m * V(1,2) +  240.560m : 
+ (V(1,2) <    5.700 ) ?    1.800m * V(1,2) +  240.560m : 
+ (V(1,2) <    5.800 ) ?    1.900m * V(1,2) +  239.990m : 
+ (V(1,2) <    5.900 ) ?    4.100m * V(1,2) +  227.230m : 
+ (V(1,2) <    6.000 ) ?   28.000m * V(1,2) +   86.220m : 
+ (V(1,2) <    6.100 ) ? -111.900m * V(1,2) +  925.620m : 
+ (V(1,2) <    6.200 ) ?   63.300m * V(1,2) + -143.100m : 
+ (V(1,2) <    6.300 ) ?   17.300m * V(1,2) +  142.100m : 
+ (V(1,2) <    6.400 ) ?    6.300m * V(1,2) +  211.400m : 
+ (V(1,2) <    6.500 ) ?    3.800m * V(1,2) +  227.400m : 
+ (V(1,2) <    7.000 ) ?    2.000m * V(1,2) +  239.100m : 
+ (V(1,2) <    7.500 ) ?    1.860m * V(1,2) +  240.080m : 
+ (V(1,2) <    8.000 ) ?    1.800m * V(1,2) +  240.530m : 
+ (V(1,2) <    8.500 ) ?    1.780m * V(1,2) +  240.690m : 
+ (V(1,2) <    9.000 ) ?    1.800m * V(1,2) +  240.520m : 
+ (V(1,2) <    9.500 ) ?    1.780m * V(1,2) +  240.700m : 
+ (V(1,2) <   10.000 ) ?    1.760m * V(1,2) +  240.890m : 
+    1.000n * V(1,2) +  258.490m
.ENDS


.SUBCKT	PWR_CLAMP	3    4   1   2
; connections:      Out+ Out In+ In
B1	3 4	I=
+ (V(1,2) <   -5.000 ) ?    1.000n * V(1,2) +   25.120  : 
+ (V(1,2) <   -4.800 ) ?   -6.150  * V(1,2) +   -5.630  : 
+ (V(1,2) <   -4.600 ) ?   -6.150  * V(1,2) +   -5.630  : 
+ (V(1,2) <   -4.400 ) ?   -6.150  * V(1,2) +   -5.630  : 
+ (V(1,2) <   -4.200 ) ?   -6.100  * V(1,2) +   -5.410  : 
+ (V(1,2) <   -4.000 ) ?   -6.150  * V(1,2) +   -5.620  : 
+ (V(1,2) <   -3.800 ) ?   -6.100  * V(1,2) +   -5.420  : 
+ (V(1,2) <   -3.600 ) ?   -6.150  * V(1,2) +   -5.610  : 
+ (V(1,2) <   -3.400 ) ?   -6.100  * V(1,2) +   -5.430  : 
+ (V(1,2) <   -3.200 ) ?   -6.150  * V(1,2) +   -5.600  : 
+ (V(1,2) <   -3.000 ) ?   -6.100  * V(1,2) +   -5.440  : 
+ (V(1,2) <   -2.800 ) ?   -6.100  * V(1,2) +   -5.440  : 
+ (V(1,2) <   -2.600 ) ?   -6.100  * V(1,2) +   -5.440  : 
+ (V(1,2) <   -2.400 ) ?   -6.100  * V(1,2) +   -5.440  : 
+ (V(1,2) <   -2.200 ) ?   -6.050  * V(1,2) +   -5.320  : 
+ (V(1,2) <   -2.000 ) ?   -6.050  * V(1,2) +   -5.320  : 
+ (V(1,2) <   -1.950 ) ?   -6.000  * V(1,2) +   -5.220  : 
+ (V(1,2) <   -1.900 ) ?   -6.200  * V(1,2) +   -5.610  : 
+ (V(1,2) <   -1.850 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.800 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.750 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.700 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.650 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.600 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.550 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.500 ) ?   -6.000  * V(1,2) +   -5.230  : 
+ (V(1,2) <   -1.450 ) ?   -5.800  * V(1,2) +   -4.930  : 
+ (V(1,2) <   -1.400 ) ?   -6.000  * V(1,2) +   -5.220  : 
+ (V(1,2) <   -1.350 ) ?   -5.800  * V(1,2) +   -4.940  : 
+ (V(1,2) <   -1.300 ) ?   -6.000  * V(1,2) +   -5.210  : 
+ (V(1,2) <   -1.250 ) ?   -5.800  * V(1,2) +   -4.950  : 
+ (V(1,2) <   -1.200 ) ?   -5.800  * V(1,2) +   -4.950  : 
+ (V(1,2) <   -1.150 ) ?   -5.600  * V(1,2) +   -4.710  : 
+ (V(1,2) <   -1.100 ) ?   -5.800  * V(1,2) +   -4.940  : 
+ (V(1,2) <   -1.050 ) ?   -5.400  * V(1,2) +   -4.500  : 
+ (V(1,2) <   -1.000 ) ?   -5.490  * V(1,2) +   -4.594  : 
+ (V(1,2) < -950.000m) ?   -4.991  * V(1,2) +   -4.096  : 
+ (V(1,2) < -900.000m) ?   -4.992  * V(1,2) +   -4.096  : 
+ (V(1,2) < -850.000m) ?   -3.383  * V(1,2) +   -2.649  : 
+ (V(1,2) < -800.000m) ?   -3.383  * V(1,2) +   -2.649  : 
+ (V(1,2) < -750.000m) ? -568.000m * V(1,2) + -396.370m : 
+ (V(1,2) < -700.000m) ? -568.200m * V(1,2) + -396.520m : 
+ (V(1,2) < -650.000m) ?  -11.990m * V(1,2) +   -7.173m : 
+ (V(1,2) < -600.000m) ?  -12.056m * V(1,2) +   -7.216m : 
+ (V(1,2) < -550.000m) ? -174.000u * V(1,2) +  -86.740u : 
+ (V(1,2) < -500.000m) ? -174.153u * V(1,2) +  -86.824u : 
+ (V(1,2) < -450.000m) ?   -2.488u * V(1,2) + -991.660n : 
+ (V(1,2) < -400.000m) ?   -2.488u * V(1,2) + -991.750n : 
+ (V(1,2) < -350.000m) ?  -36.000n * V(1,2) +  -10.870n : 
+ (V(1,2) < -300.000m) ?  -35.845n * V(1,2) +  -10.816n : 
+ (V(1,2) < -250.000m) ?  -96.400p * V(1,2) +  -91.180p : 
+ (V(1,2) < -200.000m) ?  -96.600p * V(1,2) +  -91.230p : 
+ (V(1,2) < -150.000m) ? -363.800p * V(1,2) + -144.670p : 
+ (V(1,2) < -100.000m) ? -363.800p * V(1,2) + -144.670p : 
+ (V(1,2) <  -50.000m) ?  415.800p * V(1,2) +  -66.710p : 
+ (V(1,2) <    0.000 ) ?  416.000p * V(1,2) +  -66.700p : 
+    1.000n * V(1,2) +  -66.700p
.ENDS

  
.END 
